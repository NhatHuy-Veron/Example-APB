package apb_pkg;

`include "uvm_macros.svh"
import uvm_pkg::*;

// Include all TB components
`include "apb_transaction.sv"
`include "apb_sequencer.sv"
`include "apb_driver.sv"
`include "apb_monitor.sv"
`include "apb_agent.sv"
`include "apb_environment.sv"

endpackage